module Decode(
              input clk,
              input rst
);

   always_comb begin
   end
endmodule
